`default_nettype none //do not allow undeclared wires

module risk_alu(reg1,reg2)

endmodule
module cpu(
    input wire clk,
    output wire [3:0] led
);

endmodule
